---------------------------------down-------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:22:44 02/13/2017 
-- Design Name: 
-- Module Name:    CGROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNIMACRO;
use UNIMACRO.Vcomponents.ALL;

	
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CGROM2 is


Port (

	CGROM_CLK 		: in STD_LOGIC;
	CGROM_EN 		: in STD_LOGIC;
	CGROM_ADDR 		: in STD_LOGIC_VECTOR(13 downto 0); -- change this to (11 downto 0) once we have a full character set
	CGROM_DO 		: out STD_LOGIC_VECTOR(0 downto 0);
	
	DI					: in STD_LOGIC_VECTOR(0 downto 0);
	REGCE				: in STD_LOGIC;
	RST				: in STD_LOGIC;
	WE					: in STD_LOGIC_VECTOR(0 downto 0);
	WRADDR			: in STD_LOGIC_VECTOR(13 downto 0);
	WRCLK				: in STD_LOGIC;
	WREN				: in STD_LOGIC
	);

end CGROM;

architecture Behavioral of CGROM2 is

begin
BRAM_SDP_MACRO_inst: BRAM_SDP_MACRO
generic map (
	BRAM_SIZE=>"18Kb",
	DEVICE=>"SPARTAN6",
	WRITE_WIDTH=>1,
	READ_WIDTH=>1,
	DO_REG=>0,
	INIT_FILE=>"NONE",
	SIM_COLLISION_CHECK=>"ALL",
	SIM_MODE=>"SAFE",
	SRVAL=>X"00000000000000000",
	INIT=>X"00000000000000000",

--
-- here's our ASCII 8x8 CGROM. The 3 MSBs control the scan line. 
-- right now the upper 128 characters are inverse video.
--
--
-- this is a codepage 437 font 

INIT_00=> X"000000000000181818007CFE6618400199FEFC3CF0FF00FF00081C08367E7E00", -- 00
INIT_01=> X"1E06001800001E1E3F1C3F381E1E0C3E6000000000000618061C000C36360C00",
INIT_02=> X"00081E031E7F33636333333F1E3F1E3F1C63630F67781E333C7F7F1F3C3F0C3E",
INIT_03=> X"006E07183800000000000008000000000000000E07300C07001C00380007000C",
INIT_04=> X"701F331C1833C300001E00001E7C00380C63073E3307337E000C07337E38001E",
INIT_05=> X"00186C6C006C6C00006C181818DBAA44000018C3C300000C1C3C3F0000001C38",
INIT_06=> X"FFF00F00FF0018186C0000186C00006C186C006C006C006C6C18180018001818",
INIT_07=> X"00000E1EF000001C000C187018060C001E1C6000381C1C3F0000003F00000000",
INIT_08=> X"FF1824000C18183C3C00C6DB663C70075AC6CC66E0C33CFF00083E1C7FFF8100", -- 01
INIT_09=> X"330C000C0C0C33333306033C33330E63300000000C660C0C0636633E36361E00",
INIT_0A=> X"001C1806066333636333332D336633663667770666300C336646463666661E63",
INIT_0B=> X"083B0C180C0000000000000C000000000000000C06000006003600300006000C",
INIT_0C=> X"D83333361800183307330733333600000C1C0063000000C3000C0000C3003333",
INIT_0D=> X"00186C6C006C6C00006C181818EE551133CC1863630000003636001F38380000",
INIT_0E=> X"FFF00F00FF0018186C0000186C00006C186C006C006C006C6C18180018001818",
INIT_0F=> X"00001836300000366E0C18D80C0C0C3F330630000C36360C6E6600337F3F1E00",
INIT_10=> X"FF3C66030630187E7E001CDB667E7C1F3CFEFC66F09966E7181C1C3E7FDBA500", -- 02
INIT_11=> X"30183F060C0C333330031F3630300C73180000000C3C1806031C33037F361E00",
INIT_12=> X"0036180C063133366333330C07663366636F7F0636300C33031616660366337B",
INIT_13=> X"1C000C180C3F33636333333E3E3B6E3B1E1F330C66300E366E061E301E061E18",
INIT_14=> X"18331E267E333C00000000000033FE3F00360E1C0E1E1E3C1E1E1E1E3C1E0003",
INIT_15=> X"001F6C6F7F6C6F1F006C1F1818DBAA44666600333300000C3636330000000E1E",
INIT_16=> X"FFF00F00FF0018FF6C00F8F86C00FF6CFFEFFFECFFEFFCEC6CF8180018001818",
INIT_17=> X"003C0C36300000363B0018D806183F0033037E7E1863631E3B667E063633336E",
INIT_18=> X"7E7EFF037F7F1818180036DE66187F7FE7C60C66BEBD42C33C3E7F7F7FFF8100", -- 03
INIT_19=> X"1830000300003E1E181F30331C1C0C7B0C003F003FFF1806006E181E36000C00",
INIT_1A=> X"0063181806181E1C6B33330C0E3E333E637B7F061E300C3F031E1E66033E337B",
INIT_1B=> X"36003800071933366B33330C036E336633337F0C36300C6E330F333E333E3000",
INIT_1C=> X"3C5F3F0F0333663333331E1E1E7F30061E630C180C3333660330303060333333",
INIT_1D=> X"00186C60606C6018006C181818775511CC3318DB7B3F3F061C7C371F331E0C30",
INIT_1E=> X"FFF00F00FF0018186C0018186C00006C0000000C00000C0C6C18180018001818",
INIT_1F=> X"003C06363000181C003F18180C0C0C3F331FDBDB3E637F3318661B0C36031F3B",
INIT_20=> X"3CFF660306307E187E7E36D866187C1FE7C60C3C33BD42C33C7F7F3E3EC3BD00", -- 04
INIT_21=> X"0C180006000030330C33307F30060C6F060000000C3C1806003B0C307F000C00",
INIT_22=> X"00001830064C0C1C7F33330C38363B0663736B4636330C337316166603663F7B",
INIT_23=> X"63000C180C0C331C7F33330C1E66336633337F0C1E300C6633063F3303663E00",
INIT_24=> X"18630C0603336633333333333333FE1E337F0C180C3F3F7E033E3E3E7C3F331E",
INIT_25=> X"1F1F7F7F6F6C6F1F7F6F1F1F18DBAA44666618ECCC30030300003F3333330C3E",
INIT_26=> X"00F00FFFFFF81FFFFFFCF8F8FCFFFFFFFFEFFFECEFFFECFCECF8FFFFF8FFFFF8",
INIT_27=> X"003C1E36371818006E00181818060C003303DBDB3336633318661B0636033313",
INIT_28=> X"18FF247F0C183C183C7E1CD8007E70073CE60E18339966E7183E3E1C1CE79900", -- 05
INIT_29=> X"000C3F0C0C0C18330C33333033330C67030C000C0C660C0C0033661F36000000",
INIT_2A=> X"0000186006660C36771E330C33661E063663636666330C336606463666663303",
INIT_2B=> X"63000C180C263E367F1E332C30063E3E33336B0C36330C663E06033333663300",
INIT_2C=> X"18F33F677E333C3E33333333333333063F630C180C0303061E33333366033318",
INIT_2D=> X"180000006C6C6C186C6C181818EE551133CC18F6663003333E7E3B3333330C33",
INIT_2E=> X"00F00FFFFF1800186C6C1800006C1800006C006C6C006C006C18180018180000",
INIT_2F=> X"003C0000360000003B0C1B180000003F33067E7E3336361E183E1B3336031F3B",
INIT_30=> X"0000000000001818187E33D8663C40015A670F7E33C33CFF001C1C0808FF8100", -- 06
INIT_31=> X"0C0600180C0C0E1E0C1E1E781E3F3F3E010C000C00000618006E630C36000C00",
INIT_32=> X"00001E401E7F1E63630C3F1E1E67380F1C63637F671E1E337C0F7F1F3C3F331E",
INIT_33=> X"7F000718383F3063360C6E181F0F30061E33631E67331E67300F1E6E1E3B6E00",
INIT_34=> X"1B630C3F181E18307E7E1E1E1E73FE3F33631E3C1E1E1E3C307E7E7EFC1E7E30",
INIT_35=> X"180000006C6C6C186C6C181818DBAA44000018F33300001E000033337E1E1E7E",
INIT_36=> X"00F00FFFFF1800186C6C1800006C1800006C006C6C006C006C18180018180000",
INIT_37=> X"000000003C000000000C1B183F3F3F00331C06001E771C0C18060E3F3603036E",
INIT_38=> X"0000000000000000FF001E0000180000990307181EFF00FF003E3E00007E7E00", -- 07
INIT_39=> X"0000000006000000000000000000000000000006000000000000000000000000",
INIT_3A=> X"FF00000000000000000000000000000000000000000000000000000000000000",
INIT_3B=> X"0000000000001F00000000000000780F00000000001E00001F00000000000000",
INIT_3C=> X"0EE30C001800001F000000000000000000000000000000001C0000000000001E",
INIT_3D=> X"180000006C6C6C186C6C181818775511000000C0F00000000000000000000000",
INIT_3E=> X"00F00FFFFF1800186C6C1800006C1800006C006C6C006C006C18180018180000",
INIT_3F=> X"000000003800000000000E1800000000000003000000003F0003000000000300")

--INITP_00=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_01=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_02=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_03=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_04=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_05=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_06=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_07=> X"0000000000000000000000000000000000000000000000000000000000000000")
		
	port map (
		DO=>CGROM_DO,
		DI=>DI,
		RDADDR=>CGROM_ADDR,
		RDCLK=>CGROM_CLK,
		RDEN=>CGROM_EN,
		REGCE=>REGCE,
		RST=>RST,
		WE=>WE,
		WRADDR=>WRADDR,
		WRCLK=>WRCLK,
		WREN=>WREN
		);


end Behavioral;

