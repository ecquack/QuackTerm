---------------------------------down-------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:22:44 02/13/2017 
-- Design Name: 
-- Module Name:    CGROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNIMACRO;
use UNIMACRO.Vcomponents.ALL;

	
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CGROM is


Port (

	CGROM_CLK 		: in STD_LOGIC;
	CGROM_EN 		: in STD_LOGIC;
	CGROM_ADDR 		: in STD_LOGIC_VECTOR(13 downto 0); -- change this to (11 downto 0) once we have a full character set
	CGROM_DO 		: out STD_LOGIC_VECTOR(0 downto 0);
	
	DI					: in STD_LOGIC_VECTOR(0 downto 0);
	REGCE				: in STD_LOGIC;
	RST				: in STD_LOGIC;
	WE					: in STD_LOGIC_VECTOR(0 downto 0);
	WRADDR			: in STD_LOGIC_VECTOR(13 downto 0);
	WRCLK				: in STD_LOGIC;
	WREN				: in STD_LOGIC
	);

end CGROM;

architecture Behavioral of CGROM is

begin
BRAM_SDP_MACRO_inst: BRAM_SDP_MACRO
generic map (
	BRAM_SIZE=>"18Kb",
	DEVICE=>"SPARTAN6",
	WRITE_WIDTH=>1,
	READ_WIDTH=>1,
	DO_REG=>0,
	INIT_FILE=>"NONE",
	SIM_COLLISION_CHECK=>"ALL",
	SIM_MODE=>"SAFE",
	SRVAL=>X"00000000000000000",
	INIT=>X"00000000000000000",

--
-- here's our ASCII 8x8 CGROM. The 3 MSBs control the scan line. 
-- right now the upper 128 characters are inverse video.
--
--
-- this is a codepage 850 font with out the need for the NOT in the VGA pixel calculation

--
INIT_00=> X"000000000000181818007CFE6618400118FEFC3CF0FF00FF00081C08367E7E00", -- 00
INIT_01=> X"3E06006000003E3E7F1C7F383E3E181C6000000000000C30181C001836661800",
INIT_02=> X"00083C033C7F66636363637E3C3F3E3F3E63630F67783C633C7F7F1F3C3F1C3E",
INIT_03=> X"006E0E18700000000000000C000000000000001C07601807003C00380007000C",
INIT_04=> X"70005C1C00636363061E0C633E7C00181C630C3E660C633E000C0C633E30333E",
INIT_05=> X"0066186C006C6C7E183E0C1818EEAA44000018C6C6007E181C3C6E6E18303018",
INIT_06=> X"FF0C1800FF0018663C30000C633E1F0C006C006C006C006C6E6E180018001818",
INIT_07=> X"00001E1E1800001C00007CFE8700180030FF3018063E180F07006E6E303E1E0C",
INIT_08=> X"FF1824000C18183C3C0086DB663C7007DBC6CC66E0C33CFF001C3E1C7FFF8100", -- 01
INIT_09=> X"630C0030181863636306033C63631C3630000000186618181836637C36663C00",
INIT_0A=> X"001C30060C6366636363637E6666636663677706663018636646463666663663",
INIT_0B=> X"083B1818180000000000000C0000000000000018060000060066003000060018",
INIT_0C=> X"D863363640001C000C2118004136000C361C184100180041000C180041180063",
INIT_0D=> X"0066186C006C6C813041061818BB551133CC00676700810036363B3B0C18180C",
INIT_0E=> X"FF181800FF001800421800180041367E636C006C006C006C3B3B180018001818",
INIT_0F=> X"000030301C006336001886DB4C0018001800180C0C410C0606003B3B60413306",
INIT_10=> X"FF3C66030630187E7E003CDB667E7C1F3CFEFC66F09966E7183E1C3E7FDBA500", -- 02
INIT_11=> X"30187E1818186363300303366060186318000000183C300C0C1C33067F243C00",
INIT_12=> X"0036300C0C3166366363635A0C666366636F7F0636301863031616660366637B",
INIT_13=> X"1C001818187E63636363333F7E3B6E3B3E3B371866601C366E063E3E3E3E1E30",
INIT_14=> X"183673263E63366333003E3E3E337E7F3E36001C1C3E3E3E7E1E1E1E1E3E3303",
INIT_15=> X"003C7E6F7F6C6FB91C1C1C1818EEAA446666183636009D1836360000333E001E",
INIT_16=> X"FF3C1800FF00183C3C3C1C7F7F7F66303EEFFFECFFEFFCEC1C3E180018001818",
INIT_17=> X"003C181C1800003600003CDB27007E000C0066636300633E3E661C3E1C1C331C",
INIT_18=> X"7E7EFF037F7F1818180066DE66187F7FE7C60C66BEBD42C33C7F7F7F7FFF8100", -- 03
INIT_19=> X"1830000C00007E3E183F3F333C38186B0C007E007EFF300C006E183C36001800",
INIT_1A=> X"006330180C183C1C6B636318183E633E637B7F061E30187F031E1E66033E7F7B",
INIT_1B=> X"360070180E3263366B63330C036E336663667F183660186E331F633363663000",
INIT_1C=> X"3C1C6B0F7363636333336363637F480363631C18186363630330303030633303",
INIT_1D=> X"007E0360606C60853636361818BB5511CC33185E7E7FA5181C7C673B33631C30",
INIT_1E=> X"FF180000FF0018181818180303036F3E6300000C00000C0C3660180018001818",
INIT_1F=> X"003C0C301818001C007E66DE5C00187E00006663636363666666366336361B36",
INIT_20=> X"3CFF660306307E187E7E66D866187C1FE7C60C3C33BD42C33C7F7F3E3EC3BD00", -- 04
INIT_21=> X"18180018000060630C63607F600C186306000000183C300C003B0C607F001800",
INIT_22=> X"000030300C4C18366B6363183036630663736B4636331863731616660366637B",
INIT_23=> X"630018181818631C6B63330C3E06336663666B181E60186633067F3303663E00",
INIT_24=> X"183667066B6363633333636363337F1F7F7F1818187F7F7F033E3E3E3E7F3363",
INIT_25=> X"1F18037F6F6C6F856363631F18EEAA4466663C6CCC609D0C00006F663363183E",
INIT_26=> X"001800FFFFF81F181818183F3F3F663363EFFFECEFFFECFC637EFFFFF8FFFFF8",
INIT_27=> X"003C3E1E3C000000000066D86F00180000003C636363633E6666636363633363",
INIT_28=> X"18FF247F0C183C183C7E3CD8007E70073CE60E18339966E7183E6B1C1CE79900", -- 05
INIT_29=> X"000C7E30181830630C6363306366183603180018186618180033663E36000000",
INIT_2A=> X"000030600C6618637F3663186666730663636366663318636606463666666303",
INIT_2B=> X"63001818184C7E367F36336C60063E3E63666B18366618663E06033363663300",
INIT_2C=> X"1B6336666763367E333363636333090363631818180303037E3333333303333E",
INIT_2D=> X"187E7E006C6C6CB97F7F7F1818BB551133CC3C566660A5C63E7E7B6633631833",
INIT_2E=> X"001818FFFF18001818181803030336333E6C006C6C006C007F63180018180000",
INIT_2F=> X"003C00000000000018183CD854FF00000000187E636363063E66366336366336",
INIT_30=> X"0000000000001818187E61D8663C4001DB670F7E33C33CFF0008080808FF8100", -- 06
INIT_31=> X"1806006018181E3E0C3E3E783E7F7E1C0118001800000C30006E631836001800",
INIT_32=> X"00003C403C7F3C63361C3E3C3C673E0F3E63637F671E3C635C0F7F1F3C3F631E",
INIT_33=> X"7F000E18707E6063361C6E383F0F30063E666B3C67663C67300F3E6E3E3B6E00",
INIT_34=> X"0E001D3F3E3E1C606E6E3E3E3E737F7F63633C3C3C3E3E3E306E6E6E6E3E6E30",
INIT_35=> X"181818006C6C6C816363631818EEAA44000018FB3300817C000073666E3E3C6E",
INIT_36=> X"003C18FFFF18003C3C3C3C7F7F7F1F1E636C006C6C006C00637E180018180000",
INIT_37=> X"0000000000000000300061D8FA007E0000003C603E3E3E0F063E1C3E1C1C331C",
INIT_38=> X"0000000000000000FF003E0000180000180307181EFF00FF001C1C00007E7E00", -- 07
INIT_39=> X"000000000C00000000000000000000000000000C000000000000000000000000",
INIT_3A=> X"FF00000000000000000000000000700000000000000000000000000000000000",
INIT_3B=> X"0000000000003F00000000000000780F00000000003C00001F00000000000000",
INIT_3C=> X"000000000100003F000000000000000000000000000000001C0000000000001E",
INIT_3D=> X"181818006C6C6C7E0000001818BB551100000060F0007E000000000000000000",
INIT_3E=> X"000018FFFF1800000000000000000000006C006C6C006C000000180018180000",
INIT_3F=> X"00000000000000001C003E0061FF00000000003F000000000F03000000000000")

--INITP_00=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_01=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_02=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_03=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_04=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_05=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_06=> X"0000000000000000000000000000000000000000000000000000000000000000",
--	INITP_07=> X"0000000000000000000000000000000000000000000000000000000000000000")
		
	port map (
		DO=>CGROM_DO,
		DI=>DI,
		RDADDR=>CGROM_ADDR,
		RDCLK=>CGROM_CLK,
		RDEN=>CGROM_EN,
		REGCE=>REGCE,
		RST=>RST,
		WE=>WE,
		WRADDR=>WRADDR,
		WRCLK=>WRCLK,
		WREN=>WREN
		);


end Behavioral;

